package decode_test_pkg;

	import uvm_pkg::*;
	import uvmf_base_pkg_hdl::*;
	import uvmf_base_pkg::*;
	`include "uvm_macros.svh"
	import decode_in_pkg::*;
	import decode_out_pkg::*;
	import decode_env_pkg::*;
	
	`include "src/decode_test.svh"

endpackage
